/* Definition of the `ping` component. */

component mqtt_subscriber.Ping

endpoints {
    /* Declaration of a named implementation of the "Ping" interface. */
    ping : mqtt_subscriber.Ping
}
